module top (
    input clk_25mhz
);

endmodule
