module top (
    input clk_25mhz,

    output h_sync,
    output v_sync,


    output [3:0] r,
    output [3:0] g,
    output [3:0] b
);

    

endmodule
