module Raytracer(
	input wire pixel_clk,
	input reg [10:0] x,
	input reg [10:0] y,
	output reg [2:0] rgb
);

endmodule
